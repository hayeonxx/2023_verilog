module cla(
    input [3:0] a,
    input [3:0] b,
    output c_in,
    output [3:0] s,
    output c_out
);

endmodule