module encoder(
    input alu_done,
    input [31:0] cal_result,
    output [7:0] uart_out,
    output uartout_valid
);

endmodule