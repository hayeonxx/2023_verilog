module decoder(
    input [7:0] data_out;
    input dataout_valid;
    output [3:0] data_type;
    output [1:0] op;
    output [3:0] a;
    output [3:0] b;
    output paser_done;
);



endmodule