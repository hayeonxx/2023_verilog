module testbench;

endmodule