module add(a,b,o_add);

input [15:0] a, b;
output [15:0] o_add;
assign o_add = a + b;

endmodule